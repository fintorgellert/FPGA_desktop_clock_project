`timescale 1ns / 1ps

module hexled(
    input [5:0] val,
    input rst,
    output [5:0] led
); 

    reg [5:0] disp;

    always @(*) 
        begin
            if (rst)
                disp <= 6'b0;   
            else
                disp <= val;       
        end
    
    assign led = disp;    
        
endmodule

